module vvk
